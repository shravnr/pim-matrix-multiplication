package types;

    parameter int MATRIX_SIZE = 8;
    parameter int CHUNK_SIZE = MATRIX_SIZE/2;

    parameter int LEN = 32; // Adress width
    parameter int WIDTH = 32; // Data width
    parameter int MEM_ELEMENTS = 1024;

endpackage




