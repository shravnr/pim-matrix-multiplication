module memory
import types::*;
(
    input         clk,
    input         rst,
    input logic [LEN-1:0] src1_addr,
    input logic [LEN-1:0] src2_addr,
    input logic [LEN-1:0] dst_addr,
    // input logic [2:0]     matrix_size,

    input logic start
);

    // Memory
    logic [WIDTH-1:0] mem[MEM_ELEMENTS-1:0];

    //Inputs to PIM-C
    logic [WIDTH-1:0] matrix_A [MATRIX_SIZE**2-1:0];
    logic [WIDTH-1:0] matrix_B [MATRIX_SIZE**2-1:0];
    logic [WIDTH-1:0] result [MATRIX_SIZE**2-1:0];
    logic pim_unit_start;

    //Output from PIM-C
    logic result_ready;

    //Memory FSM States
    typedef enum logic [1:0] {
        IDLE,
        READ_MATRICES,
        COMPUTE,
        WRITE_RESULT
    } state_t;

    state_t current_state, next_state;
    


    //Drive State Machine
    always_ff @(posedge clk) begin
        if(rst) current_state <= IDLE;
        else    current_state <= next_state;
    end

    //State Transition Logic
    always_comb begin
        next_state = current_state;
        case(current_state) 
            IDLE:               if(start) next_state = READ_MATRICES;
            READ_MATRICES:      next_state = COMPUTE;
            COMPUTE:            if(result_ready) next_state = WRITE_RESULT;
            WRITE_RESULT:       next_state= IDLE;
        endcase
    end

    pim_controller pim_ctl (
        .clk(clk), //clock synchronization ensured. so I don't think modules need to be called within an always_ff (i don't think that's valid either)
        .rst(rst),
        .start(pim_unit_start), 
        .matrix_A(matrix_A), 
        .matrix_B(matrix_B), 
        // .matrix_size(matrix_size),
        //.no_of_pims(no_of_pims),
        .result(result),
        .result_ready(result_ready)//output from PIM-C-- but does it need to communicate with memory? might need another wrapper here 
    );

    //State Logic
    always_ff @(posedge clk) begin
        if(rst) begin
            //DENSE
            // X X
            // X X
            for (int i = 0; i < MEM_ELEMENTS; i++) begin
                mem[i] <= i;
            end
            //SPARSE
            // one diagonal matrix from 0 
            /*
            for (int i = 0; i < MATRIX_SIZE**2; i++) begin
                automatic int row = i / MATRIX_SIZE;
                automatic int col = i % MATRIX_SIZE;
                if (row != col) begin
                    mem[i] <= 0;
                end
            end*/
            

            
            /*
            // 0 X
            // 0 X
            mem[100]<=0;
            mem[101]<=0;
            mem[104]<=0;
            mem[105]<=0;
            mem[108]<=0;
            mem[109]<=0;
            mem[112]<=0;
            mem[113]<=0;
            /*
            // X 0
            // X 0
            mem[102]<=0;
            mem[103]<=0;
            mem[106]<=0;
            mem[107]<=0;
            mem[110]<=0;
            mem[111]<=0;
            mem[114]<=0;
            mem[115]<=0; */

            /*
            //  X 0
            //  0 X
            mem[102]<=0;
            mem[103]<=0;
            mem[106]<=0;
            mem[107]<=0;
            mem[108]<=0;
            mem[109]<=0;
            mem[112]<=0;
            mem[113]<=0;
           */

            /*
            //  0 X
            //  X 0
            mem[100]<=0;
            mem[101]<=0;
            mem[104]<=0;
            mem[105]<=0;
            mem[110]<=0;
            mem[111]<=0;
            mem[114]<=0;
            mem[115]<=0;
           */

        end else begin
            case(current_state)

                IDLE: begin
                    // busy<=0;
                    // done<=0;
                end

                READ_MATRICES: begin
                    $display("Start time [%0t]", $time);

                    for (int i = 0; i < MATRIX_SIZE**2; i++) begin
                        matrix_A[i] <= mem[src1_addr + i];
                        matrix_B[i] <= mem[src2_addr + i];
                    end

                    // busy<=1;
                    pim_unit_start <= 1'b1;

                end

                COMPUTE: begin
                    pim_unit_start <= 1'b0;
                end

                WRITE_RESULT: begin

                    for (int i = 0; i < MATRIX_SIZE**2; i++) begin
                        mem[dst_addr + i] <= result[i];
                    end
                    
                    $display("End time [%0t]", $time);
                    // done<=1;
                    // busy<=0;
                end
                

            endcase
        end

    end


endmodule