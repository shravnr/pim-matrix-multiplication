package types;



endpackage




